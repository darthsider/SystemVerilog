library verilog;
use verilog.vl_types.all;
entity counter_tb_top is
end counter_tb_top;
