`include "transaction.sv"
`include "generator.sv"
`include "intf.sv"
`include "driver.sv"
`include "environment.sv"
`include "test.sv"
`include "mux.v"
`include "tbench_top.sv"

