`include "counter.v"
`include "counter_trans.sv"
`include "counter_gen.sv"
`include "counter_intf.sv"
`include "counter_bfm.sv"
`include "counter_env.sv"
`include "counter_test.sv"
`include "tb_counter_top.sv"
