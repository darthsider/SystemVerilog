library verilog;
use verilog.vl_types.all;
entity counter_test is
end counter_test;
