library verilog;
use verilog.vl_types.all;
entity comp_files_sv_unit is
end comp_files_sv_unit;
