class counter_trans;
  
  rand bit load;
  rand bit [3:0] data_in;
  rand bit up_down;
  bit [3:0] data_out;
   
endclass
